library ieee;
use ieee.std_logic_1164.all;

package Pkg_find_prime_numbers_BC_Estado is
	type Estado is (
		SL01, SL03, SL03a, SL05, SL06, SL07, SL08, SL09,  
		SL10, SL11, SL12, SL13, SL14, SL15, SL16, SL18, SL19, 
		SL20, SL22, SL23, SL24, SL24a, SL25, SL26, SL26a, SL27, SL28, SL29
	);
end package;